* NGSPICE file created from Tristate_buffer.ext - technology: sky130A

.param temp=27
.param supl = 1.8V

*Including sky130 devoce models
.lib "sky130_fd_pr/models/sky130.lib.spice" tt

Vdd vdd 0 {supl}

* Top level circuit Tristate_buffer

X0 inb in gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 out enb gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 out en out1 gnd sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X3 inb in vdd vdd sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X4 out1 inb vdd vdd sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X5 out enb out1 vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X6 out1 inb gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
C0 out1 enb 0.01fF
C1 inb in 0.03fF
C2 enb vdd 0.01fF
C3 out en 0.00fF
C4 en inb 0.01fF
C5 out1 vdd 0.07fF
C6 out enb 0.05fF
C7 inb enb 0.01fF
C8 out out1 0.17fF
C9 out vdd 0.01fF
C10 out1 inb 0.12fF
C11 inb vdd 0.13fF
C12 out inb 0.01fF
C13 en enb 0.01fF
C14 in vdd 0.03fF
C15 en out1 0.01fF
C16 en gnd 0.21fF
C17 out gnd 0.18fF
C18 out1 gnd 0.46fF
C19 inb gnd 0.58fF
C20 in gnd 0.30fF
C21 enb gnd 0.36fF
C22 vdd gnd 1.79fF

* Sources
Vin in 0 pulse(0 1.8 0 60ps 60ps 0.5ns 1ns)
Ven en 0 pulse(0 1.8 0 60ps 60ps 2ns 4ns)
Venb enb 0 pulse(1.8 0 0 60ps 60ps 2ns 4ns)

.tran 0.01p 10ns

.control
run

plot en+6 enb+4 in+2 out
.endc
.end

