magic
tech sky130A
timestamp 1606209640
<< nwell >>
rect 681 16 1236 220
rect 1138 15 1236 16
<< nmos >>
rect 760 -85 775 -43
rect 903 -85 918 -43
rect 1073 -87 1128 -72
<< pmos >>
rect 760 61 775 103
rect 903 61 918 103
rect 1076 96 1131 111
<< ndiff >>
rect 1073 -36 1128 -29
rect 718 -54 760 -43
rect 718 -71 723 -54
rect 740 -71 760 -54
rect 718 -85 760 -71
rect 775 -56 818 -43
rect 775 -73 795 -56
rect 812 -73 818 -56
rect 775 -85 818 -73
rect 861 -55 903 -43
rect 861 -72 867 -55
rect 884 -72 903 -55
rect 861 -85 903 -72
rect 918 -55 961 -43
rect 918 -72 939 -55
rect 956 -72 961 -55
rect 1073 -53 1081 -36
rect 1098 -53 1128 -36
rect 1073 -72 1128 -53
rect 918 -85 961 -72
rect 1073 -104 1128 -87
rect 1073 -121 1081 -104
rect 1098 -121 1128 -104
rect 1073 -129 1128 -121
<< pdiff >>
rect 1076 148 1131 155
rect 1076 131 1084 148
rect 1101 131 1131 148
rect 1076 111 1131 131
rect 718 91 760 103
rect 718 74 724 91
rect 741 74 760 91
rect 718 61 760 74
rect 775 91 818 103
rect 775 74 796 91
rect 813 74 818 91
rect 775 61 818 74
rect 861 92 903 103
rect 861 75 866 92
rect 883 75 903 92
rect 861 61 903 75
rect 918 91 961 103
rect 918 74 939 91
rect 956 74 961 91
rect 918 61 961 74
rect 1076 79 1131 96
rect 1076 62 1084 79
rect 1101 62 1131 79
rect 1076 55 1131 62
<< ndiffc >>
rect 723 -71 740 -54
rect 795 -73 812 -56
rect 867 -72 884 -55
rect 939 -72 956 -55
rect 1081 -53 1098 -36
rect 1081 -121 1098 -104
<< pdiffc >>
rect 1084 131 1101 148
rect 724 74 741 91
rect 796 74 813 91
rect 866 75 883 92
rect 939 74 956 91
rect 1084 62 1101 79
<< psubdiff >>
rect 722 -169 751 -152
rect 769 -169 788 -152
rect 855 -169 891 -152
rect 909 -169 921 -152
<< nsubdiff >>
rect 717 167 748 184
rect 766 167 783 184
rect 850 167 888 184
rect 906 167 919 184
<< psubdiffcont >>
rect 751 -169 769 -152
rect 891 -169 909 -152
<< nsubdiffcont >>
rect 748 167 766 184
rect 888 167 906 184
<< poly >>
rect 760 103 775 116
rect 903 103 918 116
rect 1151 113 1179 121
rect 1151 111 1157 113
rect 1063 96 1076 111
rect 1131 96 1157 111
rect 1174 96 1179 113
rect 1151 87 1179 96
rect 760 15 775 61
rect 903 16 918 61
rect 722 10 775 15
rect 722 -8 731 10
rect 748 -8 775 10
rect 722 -13 775 -8
rect 870 11 918 16
rect 870 -6 878 11
rect 895 -6 918 11
rect 870 -12 918 -6
rect 760 -43 775 -13
rect 903 -43 918 -12
rect 1143 -70 1171 -61
rect 1143 -72 1149 -70
rect 760 -98 775 -85
rect 903 -98 918 -85
rect 1060 -87 1073 -72
rect 1128 -87 1149 -72
rect 1166 -87 1171 -70
rect 1143 -95 1171 -87
<< polycont >>
rect 1157 96 1174 113
rect 731 -8 748 10
rect 878 -6 895 11
rect 1149 -87 1166 -70
<< locali >>
rect 717 167 718 184
rect 736 167 748 184
rect 766 167 783 184
rect 850 167 861 184
rect 879 167 888 184
rect 906 167 919 184
rect 718 103 735 167
rect 861 103 879 167
rect 1076 148 1109 155
rect 1076 145 1084 148
rect 1027 131 1084 145
rect 1101 131 1109 148
rect 1027 128 1109 131
rect 1076 123 1109 128
rect 1151 114 1179 121
rect 1151 113 1206 114
rect 718 91 746 103
rect 718 74 724 91
rect 741 74 746 91
rect 718 61 746 74
rect 790 91 818 103
rect 790 74 796 91
rect 813 74 818 91
rect 790 61 818 74
rect 861 92 889 103
rect 861 75 866 92
rect 883 75 889 92
rect 861 61 889 75
rect 933 91 961 103
rect 933 74 939 91
rect 956 74 961 91
rect 1151 96 1157 113
rect 1174 97 1206 113
rect 1174 96 1179 97
rect 1151 87 1179 96
rect 933 61 961 74
rect 722 10 760 15
rect 722 9 731 10
rect 695 -8 731 9
rect 748 -8 760 10
rect 722 -13 760 -8
rect 801 11 818 61
rect 944 16 961 61
rect 1076 79 1109 87
rect 1076 62 1084 79
rect 1101 62 1109 79
rect 1076 55 1109 62
rect 870 11 903 16
rect 801 -6 878 11
rect 895 -6 903 11
rect 801 -43 818 -6
rect 870 -12 903 -6
rect 944 -43 961 -1
rect 1080 14 1099 55
rect 1080 -3 1126 14
rect 1080 -29 1099 -3
rect 718 -54 746 -43
rect 718 -71 723 -54
rect 740 -71 746 -54
rect 718 -85 746 -71
rect 790 -56 818 -43
rect 790 -73 795 -56
rect 812 -73 818 -56
rect 790 -85 818 -73
rect 861 -55 889 -43
rect 861 -72 867 -55
rect 884 -72 889 -55
rect 861 -85 889 -72
rect 933 -55 961 -43
rect 933 -72 939 -55
rect 956 -72 961 -55
rect 1073 -36 1106 -29
rect 1073 -53 1081 -36
rect 1098 -53 1106 -36
rect 1073 -61 1106 -53
rect 933 -85 961 -72
rect 1143 -68 1171 -61
rect 1143 -70 1198 -68
rect 724 -152 741 -85
rect 861 -152 878 -85
rect 1143 -87 1149 -70
rect 1166 -85 1198 -70
rect 1166 -87 1171 -85
rect 1143 -95 1171 -87
rect 1073 -102 1106 -97
rect 1003 -119 1008 -102
rect 1025 -104 1106 -102
rect 1025 -119 1081 -104
rect 1073 -121 1081 -119
rect 1098 -121 1106 -104
rect 1073 -129 1106 -121
rect 722 -169 724 -152
rect 741 -169 751 -152
rect 769 -169 788 -152
rect 855 -169 861 -152
rect 878 -169 891 -152
rect 909 -169 921 -152
<< viali >>
rect 718 167 736 184
rect 861 167 879 184
rect 1009 128 1027 145
rect 944 -1 961 16
rect 1008 -119 1025 -102
rect 724 -169 741 -152
rect 861 -169 878 -152
<< metal1 >>
rect 712 184 936 188
rect 712 167 718 184
rect 736 167 861 184
rect 879 167 936 184
rect 712 163 936 167
rect 1003 145 1033 151
rect 1003 128 1009 145
rect 1027 128 1033 145
rect 1003 22 1033 128
rect 937 16 1033 22
rect 937 -1 944 16
rect 961 -1 1033 16
rect 937 -7 1033 -1
rect 1003 -102 1033 -7
rect 1003 -119 1008 -102
rect 1025 -119 1033 -102
rect 1003 -125 1033 -119
rect 715 -152 931 -148
rect 715 -169 724 -152
rect 741 -169 861 -152
rect 878 -169 931 -152
rect 715 -173 931 -169
<< labels >>
flabel locali 1189 -77 1189 -77 0 FreeSans 120 0 0 0 en
flabel locali 1185 106 1185 106 0 FreeSans 120 180 0 0 enb
flabel locali 809 3 809 3 0 FreeSans 120 0 0 0 inb
flabel locali 698 0 698 0 0 FreeSans 120 0 0 0 in
flabel locali 1104 6 1104 6 0 FreeSans 120 0 0 0 out
flabel metal1 971 7 971 7 0 FreeSans 120 0 0 0 out1
flabel metal1 812 176 812 176 0 FreeSans 152 0 0 0 vdd
flabel metal1 829 -164 829 -164 0 FreeSans 152 0 0 0 gnd
<< end >>
