magic
tech sky130A
timestamp 1606021460
<< nwell >>
rect -26 141 412 180
rect -26 2 413 141
rect -26 1 366 2
<< nmos >>
rect 36 -158 51 -74
rect 174 -157 189 -73
rect 321 -116 336 -74
rect 110 -281 125 -239
<< pmos >>
rect 35 24 50 108
rect 176 23 191 107
rect 321 29 336 71
<< ndiff >>
rect -6 -130 36 -74
rect -6 -152 2 -130
rect 19 -152 36 -130
rect -6 -158 36 -152
rect 51 -80 93 -74
rect 51 -102 66 -80
rect 83 -102 93 -80
rect 51 -158 93 -102
rect 132 -129 174 -73
rect 132 -151 140 -129
rect 157 -151 174 -129
rect 132 -157 174 -151
rect 189 -129 231 -73
rect 275 -89 321 -74
rect 275 -111 283 -89
rect 300 -111 321 -89
rect 275 -116 321 -111
rect 336 -78 375 -74
rect 336 -100 351 -78
rect 368 -100 375 -78
rect 336 -116 375 -100
rect 189 -151 206 -129
rect 223 -151 231 -129
rect 189 -157 231 -151
rect 68 -253 110 -239
rect 68 -275 76 -253
rect 93 -275 110 -253
rect 68 -281 110 -275
rect 125 -245 168 -239
rect 125 -267 140 -245
rect 157 -267 168 -245
rect 125 -281 168 -267
<< pdiff >>
rect -8 63 35 108
rect -8 32 0 63
rect 18 32 35 63
rect -8 24 35 32
rect 50 62 91 108
rect 50 31 65 62
rect 83 31 91 62
rect 50 24 91 31
rect 133 62 176 107
rect 133 31 140 62
rect 158 31 176 62
rect 133 23 176 31
rect 191 62 232 107
rect 191 31 207 62
rect 225 31 232 62
rect 191 23 232 31
rect 278 63 321 71
rect 278 39 284 63
rect 301 39 321 63
rect 278 29 321 39
rect 336 63 377 71
rect 336 39 353 63
rect 370 39 377 63
rect 336 29 377 39
<< ndiffc >>
rect 2 -152 19 -130
rect 66 -102 83 -80
rect 140 -151 157 -129
rect 283 -111 300 -89
rect 351 -100 368 -78
rect 206 -151 223 -129
rect 76 -275 93 -253
rect 140 -267 157 -245
<< pdiffc >>
rect 0 32 18 63
rect 65 31 83 62
rect 140 31 158 62
rect 207 31 225 62
rect 284 39 301 63
rect 353 39 370 63
<< psubdiff >>
rect 92 -341 112 -324
rect 130 -341 249 -324
rect 266 -341 296 -324
<< nsubdiff >>
rect 0 139 37 156
rect 55 139 161 156
rect 179 139 249 156
rect 267 139 303 156
<< psubdiffcont >>
rect 112 -341 130 -324
rect 249 -341 266 -324
<< nsubdiffcont >>
rect 37 139 55 156
rect 161 139 179 156
rect 249 139 267 156
<< poly >>
rect 35 108 50 121
rect 176 107 191 121
rect 35 -5 50 24
rect 321 71 336 84
rect 176 -5 191 23
rect 35 -13 191 -5
rect 35 -20 65 -13
rect 59 -30 65 -20
rect 83 -20 191 -13
rect 265 -20 296 -10
rect 83 -30 89 -20
rect 59 -38 89 -30
rect 265 -37 271 -20
rect 289 -22 296 -20
rect 321 -22 336 29
rect 289 -37 336 -22
rect 265 -46 296 -37
rect 36 -74 51 -61
rect 174 -73 189 -60
rect 321 -74 336 -37
rect 321 -129 336 -116
rect -71 -168 -40 -158
rect 36 -168 51 -158
rect -71 -185 -63 -168
rect -45 -183 51 -168
rect 174 -182 189 -157
rect 332 -181 363 -171
rect 332 -182 339 -181
rect -45 -185 -40 -183
rect -71 -194 -40 -185
rect 174 -197 339 -182
rect 332 -198 339 -197
rect 356 -198 363 -181
rect 332 -207 363 -198
rect -10 -230 125 -215
rect -10 -251 5 -230
rect 110 -239 125 -230
rect -18 -261 13 -251
rect -18 -278 -12 -261
rect 6 -278 13 -261
rect -18 -287 13 -278
rect 110 -294 125 -281
<< polycont >>
rect 65 -30 83 -13
rect 271 -37 289 -20
rect -63 -185 -45 -168
rect 339 -198 356 -181
rect -12 -278 6 -261
<< locali >>
rect 0 139 6 156
rect 24 139 37 156
rect 55 139 137 156
rect 154 139 161 156
rect 179 139 249 156
rect 267 139 284 156
rect 0 71 17 139
rect -8 63 25 71
rect -8 32 0 63
rect 18 32 25 63
rect -8 24 25 32
rect 59 62 91 71
rect 138 70 155 139
rect 285 71 302 139
rect 59 31 65 62
rect 83 31 91 62
rect 59 24 91 31
rect 133 62 165 70
rect 133 31 140 62
rect 158 31 165 62
rect 65 -5 82 24
rect 133 23 165 31
rect 200 62 232 70
rect 200 31 207 62
rect 225 31 232 62
rect 200 23 232 31
rect 278 63 310 71
rect 278 39 284 63
rect 301 39 310 63
rect 278 29 310 39
rect 345 63 377 71
rect 345 39 353 63
rect 370 39 377 63
rect 345 29 377 39
rect 59 -13 89 -5
rect 59 -30 65 -13
rect 83 -30 89 -13
rect 59 -38 89 -30
rect 206 -24 223 23
rect 265 -20 296 -10
rect 265 -24 271 -20
rect 206 -37 271 -24
rect 289 -37 296 -20
rect 65 -74 82 -38
rect 206 -41 296 -37
rect 57 -80 93 -74
rect 57 -102 66 -80
rect 83 -102 93 -80
rect 57 -108 93 -102
rect 206 -123 223 -41
rect 265 -46 296 -41
rect 351 -20 368 29
rect 351 -37 382 -20
rect 351 -74 368 -37
rect 341 -78 375 -74
rect 275 -89 312 -82
rect 275 -111 283 -89
rect 300 -111 312 -89
rect 341 -100 351 -78
rect 368 -100 375 -78
rect 341 -108 375 -100
rect 275 -116 312 -111
rect -6 -130 30 -124
rect -6 -152 2 -130
rect 19 -152 30 -130
rect -6 -158 30 -152
rect 132 -129 168 -123
rect 132 -151 140 -129
rect 157 -151 168 -129
rect 132 -157 168 -151
rect 196 -129 231 -123
rect 196 -151 206 -129
rect 223 -151 231 -129
rect 196 -157 231 -151
rect -71 -167 -40 -158
rect -93 -168 -40 -167
rect -93 -184 -63 -168
rect -71 -185 -63 -184
rect -45 -185 -40 -168
rect -71 -194 -40 -185
rect 3 -188 20 -158
rect 140 -188 157 -157
rect 3 -205 157 -188
rect 140 -239 157 -205
rect 132 -245 168 -239
rect -18 -261 13 -251
rect -18 -278 -12 -261
rect 6 -278 13 -261
rect -18 -287 13 -278
rect 68 -253 104 -247
rect 68 -275 76 -253
rect 93 -275 104 -253
rect 132 -267 140 -245
rect 157 -267 168 -245
rect 132 -273 168 -267
rect 68 -281 104 -275
rect -10 -304 7 -287
rect 76 -324 93 -281
rect 282 -324 299 -116
rect 332 -180 363 -171
rect 332 -181 385 -180
rect 332 -198 339 -181
rect 356 -197 385 -181
rect 356 -198 363 -197
rect 332 -207 363 -198
rect 93 -341 112 -324
rect 130 -341 249 -324
rect 266 -341 282 -324
rect 278 -345 299 -341
<< viali >>
rect 6 139 24 156
rect 137 139 154 156
rect 284 139 302 156
rect 76 -341 93 -324
rect 282 -341 299 -324
<< metal1 >>
rect 0 156 308 166
rect 0 139 6 156
rect 24 139 137 156
rect 154 139 284 156
rect 302 139 308 156
rect 0 130 308 139
rect 282 -320 299 -315
rect 59 -324 305 -320
rect 59 -341 76 -324
rect 93 -341 282 -324
rect 299 -341 305 -324
rect 59 -345 305 -341
rect 278 -347 305 -345
<< labels >>
flabel metal1 62 140 110 155 0 FreeSans 152 0 0 0 vdd
flabel locali 206 -40 242 -25 0 FreeSans 120 0 0 0 dout1
flabel locali 352 -36 380 -21 0 FreeSans 104 0 0 0 dout
flabel locali 364 -196 384 -181 0 FreeSans 120 0 0 0 bl
flabel locali -92 -183 -73 -168 0 FreeSans 96 0 0 0 blbar
flabel locali -9 -303 6 -288 0 FreeSans 96 0 0 0 ren
flabel locali 66 -62 81 -44 0 FreeSans 96 0 0 0 2
flabel locali 96 -204 121 -189 0 FreeSans 96 0 0 0 3
flabel metal1 142 -340 195 -325 0 FreeSans 152 0 0 0 gnd
<< end >>
