*Model Description
.param temp=27
.param supl = 1.8V

*Including sky130 device model
.lib "sky130_fd_pr/models/sky130.lib.spice" tt

Vdd vdd 0 {supl}

* Cross-coupled transistors
XM1 q qbar vdd vdd sky130_fd_pr__pfet_01v8 w=.42 l=.15 m=1
XM2 q qbar 0 0 sky130_fd_pr__nfet_01v8 w=.84 l=.15 m=1
XM3 qbar q vdd vdd sky130_fd_pr__pfet_01v8 w=.42 l=.15 m=1
XM4 qbar q 0 0 sky130_fd_pr__nfet_01v8 w=.84 l=.15 m=1

*Access Transistors
XM5 bl wl q 0 sky130_fd_pr__nfet_01v8 w=.42 l=.15 m=1
XM6 blbar wl qbar 0 sky130_fd_pr__nfet_01v8 w=.42 l=.15 m=1

*Test Pulses
vin q 0 dc 1.8v
vwl wl 0 dc 1.8v
vbl bl 0 dc 1.8v
v2 blbar 0 dc 1.8v


.dc vin 0 1.8 0.01
.control
run 
plot -I(vin)
.endc
.end
