magic
tech sky130A
timestamp 1607217454
<< nwell >>
rect -41 -23 248 119
<< nmos >>
rect 18 -190 33 -148
rect 167 -190 182 -148
rect -27 -331 15 -316
rect 119 -331 161 -316
<< pmos >>
rect 18 -3 33 39
rect 167 -3 182 39
<< ndiff >>
rect -22 -160 18 -148
rect -22 -178 -15 -160
rect 2 -178 18 -160
rect -22 -190 18 -178
rect 33 -160 71 -148
rect 33 -178 48 -160
rect 65 -178 71 -160
rect 33 -190 71 -178
rect 127 -156 167 -148
rect 127 -179 132 -156
rect 149 -179 167 -156
rect 127 -190 167 -179
rect 182 -155 218 -148
rect 182 -178 196 -155
rect 213 -178 218 -155
rect 182 -190 218 -178
rect -27 -284 15 -278
rect -27 -301 -17 -284
rect 4 -301 15 -284
rect -27 -316 15 -301
rect 119 -283 161 -278
rect 119 -300 129 -283
rect 150 -300 161 -283
rect 119 -316 161 -300
rect -27 -348 15 -331
rect -27 -365 -18 -348
rect 3 -365 15 -348
rect 119 -345 161 -331
rect -27 -372 15 -365
rect 119 -362 128 -345
rect 149 -362 161 -345
rect 119 -371 161 -362
<< pdiff >>
rect -22 32 18 39
rect -22 4 -14 32
rect 3 4 18 32
rect -22 -3 18 4
rect 33 33 72 39
rect 33 5 47 33
rect 64 5 72 33
rect 33 -3 72 5
rect 127 30 167 39
rect 127 5 135 30
rect 152 5 167 30
rect 127 -3 167 5
rect 182 31 218 39
rect 182 6 196 31
rect 213 6 218 31
rect 182 -3 218 6
<< ndiffc >>
rect -15 -178 2 -160
rect 48 -178 65 -160
rect 132 -179 149 -156
rect 196 -178 213 -155
rect -17 -301 4 -284
rect 129 -300 150 -283
rect -18 -365 3 -348
rect 128 -362 149 -345
<< pdiffc >>
rect -14 4 3 32
rect 47 5 64 33
rect 135 5 152 30
rect 196 6 213 31
<< psubdiff >>
rect 119 -226 144 -224
rect -21 -245 21 -226
rect 44 -245 83 -226
rect 106 -245 167 -226
rect 119 -248 144 -245
<< nsubdiff >>
rect -22 70 17 94
rect 41 70 100 94
rect 124 70 190 94
<< psubdiffcont >>
rect 21 -245 44 -226
rect 83 -245 106 -226
<< nsubdiffcont >>
rect 17 70 41 94
rect 100 70 124 94
<< poly >>
rect 18 39 33 54
rect 167 39 182 54
rect 18 -38 33 -3
rect 97 -36 128 -27
rect 97 -38 104 -36
rect 18 -53 104 -38
rect 123 -53 128 -36
rect 18 -148 33 -53
rect 97 -62 128 -53
rect 95 -96 127 -88
rect 167 -96 182 -3
rect 95 -113 102 -96
rect 120 -111 182 -96
rect 120 -113 127 -111
rect 95 -121 127 -113
rect 167 -148 182 -111
rect 18 -203 33 -190
rect 167 -203 182 -190
rect -43 -331 -27 -316
rect 15 -331 119 -316
rect 161 -331 174 -316
rect 64 -358 79 -331
rect 56 -366 87 -358
rect 56 -383 63 -366
rect 81 -383 87 -366
rect 56 -391 87 -383
<< polycont >>
rect 104 -53 123 -36
rect 102 -113 120 -96
rect 63 -383 81 -366
<< locali >>
rect -26 94 190 99
rect -26 93 17 94
rect -26 69 -15 93
rect 9 70 17 93
rect 41 70 100 94
rect 124 93 190 94
rect 124 70 131 93
rect 9 69 131 70
rect 155 69 190 93
rect -26 63 190 69
rect -14 39 3 63
rect 135 39 152 63
rect -22 32 11 39
rect -22 4 -14 32
rect 3 4 11 32
rect -22 -3 11 4
rect 39 33 72 39
rect 39 5 47 33
rect 64 5 72 33
rect 39 -3 72 5
rect 127 30 160 39
rect 127 5 135 30
rect 152 5 160 30
rect 127 -3 160 5
rect 188 31 218 39
rect 188 6 196 31
rect 213 6 218 31
rect 188 -3 218 6
rect 49 -71 66 -3
rect 97 -36 128 -27
rect 196 -36 213 -3
rect 97 -53 104 -36
rect 123 -53 213 -36
rect 97 -62 128 -53
rect -72 -88 66 -71
rect -72 -286 -55 -88
rect 49 -96 66 -88
rect 95 -96 127 -88
rect 49 -113 102 -96
rect 120 -113 127 -96
rect 49 -148 66 -113
rect 95 -121 127 -113
rect 196 -148 213 -53
rect -22 -160 9 -148
rect -22 -178 -15 -160
rect 2 -178 9 -160
rect -22 -190 9 -178
rect 40 -160 71 -148
rect 40 -178 48 -160
rect 65 -178 71 -160
rect 40 -190 71 -178
rect 127 -156 158 -148
rect 127 -179 132 -156
rect 149 -179 158 -156
rect 127 -190 158 -179
rect 189 -155 218 -148
rect 189 -178 196 -155
rect 213 -178 218 -155
rect 189 -190 218 -178
rect -8 -218 9 -190
rect 133 -213 150 -190
rect 133 -218 167 -213
rect -33 -223 167 -218
rect -33 -247 -14 -223
rect 11 -224 167 -223
rect 11 -226 124 -224
rect 11 -245 21 -226
rect 44 -245 83 -226
rect 106 -245 124 -226
rect 11 -247 124 -245
rect -33 -248 124 -247
rect 149 -248 167 -224
rect -33 -252 167 -248
rect -27 -284 15 -278
rect -27 -286 -17 -284
rect -72 -301 -17 -286
rect 4 -301 15 -284
rect -72 -303 15 -301
rect -27 -308 15 -303
rect 119 -280 161 -278
rect 197 -280 214 -190
rect 119 -283 214 -280
rect 119 -300 129 -283
rect 150 -297 214 -283
rect 150 -300 161 -297
rect 119 -305 161 -300
rect -27 -348 15 -342
rect -27 -352 -18 -348
rect -54 -365 -18 -352
rect 3 -365 15 -348
rect 119 -345 161 -339
rect -54 -369 15 -365
rect -27 -372 15 -369
rect 56 -366 87 -358
rect 56 -383 63 -366
rect 81 -383 87 -366
rect 119 -362 128 -345
rect 149 -346 161 -345
rect 149 -362 193 -346
rect 119 -363 193 -362
rect 119 -371 161 -363
rect 56 -391 87 -383
rect 63 -413 81 -391
<< viali >>
rect -15 69 9 93
rect 131 69 155 93
rect -14 -247 11 -223
rect 124 -248 149 -224
<< metal1 >>
rect -32 93 190 106
rect -32 69 -15 93
rect 9 69 131 93
rect 155 69 190 93
rect -32 59 190 69
rect -33 -223 167 -213
rect -33 -247 -14 -223
rect 11 -224 167 -223
rect 11 -247 124 -224
rect -33 -248 124 -247
rect 149 -248 167 -224
rect -33 -255 167 -248
<< labels >>
flabel metal1 45 65 99 94 0 FreeSans 152 0 0 0 vdd
flabel locali 184 -51 213 -37 0 FreeSans 104 0 0 0 qbar
flabel locali -49 -87 -25 -72 0 FreeSans 104 0 0 0 q
flabel metal1 46 -243 81 -226 0 FreeSans 120 0 0 0 gnd
flabel locali 64 -407 79 -393 0 FreeSans 72 0 0 0 wl
flabel locali 168 -363 184 -346 0 FreeSans 40 0 0 0 blbar_noconn
flabel locali -53 -369 -40 -352 0 FreeSans 40 0 0 0 bl_noconn
<< end >>
