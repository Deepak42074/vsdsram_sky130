* NGSPICE file created from Tristate_buffer.ext - technology: sky130A


* Top level circuit Tristate_buffer

X0 inb in gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 out en out1 gnd sky130_fd_pr__nfet_01v8 w=550000u l=150000u
X2 inb in vdd vdd sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X3 out1 inb vdd vdd sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X4 out enb out1 vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X5 out1 inb gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
C0 out out1 0.18fF
C1 enb vdd 0.01fF
C2 in inb 0.06fF
C3 out vdd 0.01fF
C4 in out1 0.01fF
C5 en inb 0.01fF
C6 out1 inb 0.08fF
C7 en out1 0.00fF
C8 in vdd 0.03fF
C9 inb vdd 0.13fF
C10 out enb 0.00fF
C11 out1 vdd 0.08fF
C12 inb enb 0.01fF
C13 en enb 0.01fF
C14 out inb 0.01fF
C15 out1 enb 0.00fF
C16 en out 0.00fF
C17 en gnd 0.21fF
C18 out gnd 0.19fF
C19 out1 gnd 0.43fF
C20 inb gnd 0.59fF
C21 in gnd 0.30fF
C22 enb gnd 0.21fF
C23 vdd gnd 1.96fF
.end

