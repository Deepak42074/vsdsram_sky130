magic
tech sky130A
timestamp 1605954624
<< nwell >>
rect -761 38 601 226
rect -761 33 561 38
rect -761 32 2 33
rect -761 31 -133 32
rect -761 26 -134 31
rect -624 25 -481 26
<< nmos >>
rect -698 -89 -683 -47
rect -524 -90 -509 -48
rect -360 -90 -345 -48
rect -215 -90 -200 -48
rect -78 -89 -63 -47
rect 62 -89 77 -47
rect 205 -89 220 -47
rect 344 -89 359 -47
rect 481 -89 496 -47
<< pmos >>
rect -698 53 -683 108
rect -526 53 -511 108
rect -360 53 -345 108
rect -215 53 -200 108
rect -80 53 -65 108
rect 64 53 79 108
rect 205 53 220 108
rect 344 53 359 108
rect 481 53 498 108
<< ndiff >>
rect -741 -60 -698 -47
rect -741 -77 -733 -60
rect -716 -77 -698 -60
rect -741 -89 -698 -77
rect -683 -57 -640 -47
rect -683 -74 -666 -57
rect -649 -74 -640 -57
rect -683 -89 -640 -74
rect -568 -57 -524 -48
rect -568 -74 -560 -57
rect -543 -74 -524 -57
rect -568 -90 -524 -74
rect -509 -58 -464 -48
rect -509 -75 -489 -58
rect -472 -75 -464 -58
rect -509 -90 -464 -75
rect -403 -60 -360 -48
rect -403 -77 -395 -60
rect -378 -77 -360 -60
rect -403 -90 -360 -77
rect -345 -57 -299 -48
rect -345 -74 -328 -57
rect -311 -74 -299 -57
rect -345 -90 -299 -74
rect -257 -59 -215 -48
rect -257 -76 -248 -59
rect -231 -76 -215 -59
rect -257 -90 -215 -76
rect -200 -60 -153 -48
rect -200 -77 -180 -60
rect -163 -77 -153 -60
rect -200 -90 -153 -77
rect -122 -58 -78 -47
rect -122 -75 -114 -58
rect -97 -75 -78 -58
rect -122 -89 -78 -75
rect -63 -58 -18 -47
rect -63 -75 -43 -58
rect -26 -75 -18 -58
rect -63 -89 -18 -75
rect 20 -57 62 -47
rect 20 -74 27 -57
rect 44 -74 62 -57
rect 20 -89 62 -74
rect 77 -59 124 -47
rect 77 -76 100 -59
rect 117 -76 124 -59
rect 77 -89 124 -76
rect 161 -60 205 -47
rect 161 -77 170 -60
rect 187 -77 205 -60
rect 161 -89 205 -77
rect 220 -57 265 -47
rect 220 -74 237 -57
rect 254 -74 265 -57
rect 220 -89 265 -74
rect 300 -60 344 -47
rect 300 -77 309 -60
rect 326 -77 344 -60
rect 300 -89 344 -77
rect 359 -57 404 -47
rect 359 -74 376 -57
rect 393 -74 404 -57
rect 359 -89 404 -74
rect 439 -57 481 -47
rect 439 -74 446 -57
rect 463 -74 481 -57
rect 439 -89 481 -74
rect 496 -58 543 -47
rect 496 -75 519 -58
rect 536 -75 543 -58
rect 496 -89 543 -75
<< pdiff >>
rect -743 84 -698 108
rect -743 64 -735 84
rect -717 64 -698 84
rect -743 53 -698 64
rect -683 84 -639 108
rect -683 64 -663 84
rect -645 64 -639 84
rect -683 53 -639 64
rect -568 91 -526 108
rect -568 61 -561 91
rect -543 61 -526 91
rect -568 53 -526 61
rect -511 91 -464 108
rect -511 61 -490 91
rect -472 61 -464 91
rect -511 53 -464 61
rect -405 91 -360 108
rect -405 61 -398 91
rect -380 61 -360 91
rect -405 53 -360 61
rect -345 91 -301 108
rect -345 61 -328 91
rect -310 61 -301 91
rect -345 53 -301 61
rect -257 92 -215 108
rect -257 62 -249 92
rect -231 62 -215 92
rect -257 53 -215 62
rect -200 91 -153 108
rect -200 61 -179 91
rect -161 61 -153 91
rect -200 53 -153 61
rect -124 91 -80 108
rect -124 61 -117 91
rect -99 61 -80 91
rect -124 53 -80 61
rect -65 99 -20 108
rect -65 91 -18 99
rect -65 61 -44 91
rect -26 61 -18 91
rect -65 53 -18 61
rect 20 91 64 108
rect 20 61 27 91
rect 45 61 64 91
rect 20 53 64 61
rect 79 91 124 108
rect 79 61 100 91
rect 118 61 124 91
rect 79 53 124 61
rect 160 91 205 108
rect 160 61 168 91
rect 186 61 205 91
rect 160 53 205 61
rect 220 91 264 108
rect 220 61 238 91
rect 256 61 264 91
rect 220 53 264 61
rect 299 91 344 108
rect 299 61 308 91
rect 326 61 344 91
rect 299 53 344 61
rect 359 91 403 108
rect 359 61 378 91
rect 396 61 403 91
rect 359 53 403 61
rect 439 91 481 108
rect 439 61 445 91
rect 463 61 481 91
rect 439 53 481 61
rect 498 91 543 108
rect 498 61 518 91
rect 536 61 543 91
rect 498 53 543 61
<< ndiffc >>
rect -733 -77 -716 -60
rect -666 -74 -649 -57
rect -560 -74 -543 -57
rect -489 -75 -472 -58
rect -395 -77 -378 -60
rect -328 -74 -311 -57
rect -248 -76 -231 -59
rect -180 -77 -163 -60
rect -114 -75 -97 -58
rect -43 -75 -26 -58
rect 27 -74 44 -57
rect 100 -76 117 -59
rect 170 -77 187 -60
rect 237 -74 254 -57
rect 309 -77 326 -60
rect 376 -74 393 -57
rect 446 -74 463 -57
rect 519 -75 536 -58
<< pdiffc >>
rect -735 64 -717 84
rect -663 64 -645 84
rect -561 61 -543 91
rect -490 61 -472 91
rect -398 61 -380 91
rect -328 61 -310 91
rect -249 62 -231 92
rect -179 61 -161 91
rect -117 61 -99 91
rect -44 61 -26 91
rect 27 61 45 91
rect 100 61 118 91
rect 168 61 186 91
rect 238 61 256 91
rect 308 61 326 91
rect 378 61 396 91
rect 445 61 463 91
rect 518 61 536 91
<< psubdiff >>
rect -744 -167 -710 -150
rect -693 -167 -374 -150
rect -357 -167 -278 -150
rect -261 -167 196 -150
rect 213 -167 273 -150
rect 290 -167 341 -150
<< nsubdiff >>
rect -742 191 -708 208
rect -691 191 -374 208
rect -357 191 -224 208
rect -207 191 194 208
rect 211 191 333 208
rect 350 191 364 208
<< psubdiffcont >>
rect -710 -167 -693 -150
rect -374 -167 -357 -150
rect -278 -167 -261 -150
rect 196 -167 213 -150
rect 273 -167 290 -150
<< nsubdiffcont >>
rect -708 191 -691 208
rect -374 191 -357 208
rect -224 191 -207 208
rect 194 191 211 208
rect 333 191 350 208
<< poly >>
rect -216 155 -185 163
rect -216 138 -209 155
rect -192 138 -185 155
rect -698 120 -511 135
rect -216 127 -185 138
rect -698 108 -683 120
rect -526 108 -511 120
rect -360 108 -345 121
rect -215 108 -200 127
rect -80 108 -65 121
rect 64 108 79 121
rect 205 108 220 122
rect 344 108 359 121
rect 481 116 579 131
rect 481 108 498 116
rect -754 -8 -719 0
rect -754 -25 -746 -8
rect -729 -10 -719 -8
rect -698 -10 -683 53
rect -526 40 -511 53
rect -416 16 -381 24
rect -416 -1 -408 16
rect -391 14 -381 16
rect -360 14 -345 53
rect -391 -1 -345 14
rect -729 -25 -683 -10
rect -754 -31 -719 -25
rect -698 -47 -683 -25
rect -533 -11 -498 -2
rect -416 -7 -381 -1
rect -533 -28 -525 -11
rect -508 -28 -498 -11
rect -533 -35 -498 -28
rect -524 -48 -509 -35
rect -360 -48 -345 -1
rect -268 14 -237 25
rect -268 -3 -262 14
rect -245 13 -237 14
rect -215 13 -200 53
rect -80 24 -65 53
rect 64 31 79 53
rect -245 -2 -200 13
rect -245 -3 -237 -2
rect -268 -11 -237 -3
rect -215 -48 -200 -2
rect -87 16 -57 24
rect -87 -1 -81 16
rect -64 -1 -57 16
rect -87 -9 -57 -1
rect 57 23 87 31
rect 57 6 63 23
rect 80 6 87 23
rect 57 -2 87 6
rect 146 16 181 22
rect 146 -1 155 16
rect 172 14 181 16
rect 205 14 220 53
rect 172 -1 220 14
rect 146 -9 181 -1
rect -78 -47 -63 -34
rect 62 -47 77 -34
rect 205 -47 220 -1
rect 285 16 320 23
rect 285 -1 294 16
rect 311 14 320 16
rect 344 14 359 53
rect 481 40 498 53
rect 311 -1 359 14
rect 285 -8 320 -1
rect 344 -47 359 -1
rect 477 -10 507 -2
rect 477 -27 483 -10
rect 500 -27 507 -10
rect 477 -35 507 -27
rect 481 -47 496 -35
rect -698 -124 -683 -89
rect -524 -103 -509 -90
rect -360 -103 -345 -90
rect -215 -103 -200 -90
rect -78 -124 -63 -89
rect 62 -124 77 -89
rect 205 -102 220 -89
rect 344 -102 359 -89
rect 481 -102 496 -89
rect 564 -124 579 116
rect -698 -139 579 -124
<< polycont >>
rect -209 138 -192 155
rect -746 -25 -729 -8
rect -408 -1 -391 16
rect -525 -28 -508 -11
rect -262 -3 -245 14
rect -81 -1 -64 16
rect 63 6 80 23
rect 155 -1 172 16
rect 294 -1 311 16
rect 483 -27 500 -10
<< locali >>
rect -742 191 -735 208
rect -718 191 -708 208
rect -691 191 -397 208
rect -380 191 -374 208
rect -357 191 -252 208
rect -235 191 -224 208
rect -207 191 168 208
rect 185 191 194 208
rect 211 191 307 208
rect 324 191 333 208
rect 350 191 364 208
rect -735 95 -718 191
rect -397 99 -380 191
rect -252 99 -235 191
rect -216 155 -185 163
rect -216 138 -209 155
rect -192 138 -185 155
rect -216 127 -185 138
rect 20 99 37 135
rect 168 99 185 191
rect 307 99 324 191
rect -743 84 -709 95
rect -743 64 -735 84
rect -717 64 -709 84
rect -743 53 -709 64
rect -673 84 -639 95
rect -673 64 -663 84
rect -645 64 -639 84
rect -673 53 -639 64
rect -568 91 -537 99
rect -568 61 -561 91
rect -543 61 -537 91
rect -568 53 -537 61
rect -495 91 -464 99
rect -495 61 -490 91
rect -472 61 -464 91
rect -495 53 -464 61
rect -405 91 -371 99
rect -405 61 -398 91
rect -380 61 -371 91
rect -405 53 -371 61
rect -335 91 -301 99
rect -335 61 -328 91
rect -310 61 -301 91
rect -335 53 -301 61
rect -257 92 -223 99
rect -257 62 -249 92
rect -231 62 -223 92
rect -257 53 -223 62
rect -187 91 -153 99
rect -187 61 -179 91
rect -161 61 -153 91
rect -187 53 -153 61
rect -124 91 -93 99
rect -124 61 -117 91
rect -99 61 -93 91
rect -124 53 -93 61
rect -51 91 -18 99
rect -51 61 -44 91
rect -26 61 -18 91
rect -51 53 -18 61
rect -809 26 -787 43
rect -770 26 -759 43
rect -754 -8 -719 0
rect -778 -25 -746 -8
rect -729 -25 -719 -8
rect -754 -31 -719 -25
rect -667 -11 -650 53
rect -568 41 -551 53
rect -616 24 -606 41
rect -589 24 -551 41
rect -667 -28 -644 -11
rect -627 -28 -610 -11
rect -667 -52 -650 -28
rect -568 -52 -551 24
rect -481 16 -464 53
rect -416 16 -381 24
rect -481 -1 -408 16
rect -391 -1 -381 16
rect -533 -11 -498 -2
rect -533 -28 -525 -11
rect -508 -28 -498 -11
rect -533 -35 -498 -28
rect -481 -52 -464 -1
rect -416 -7 -381 -1
rect -329 15 -312 53
rect -268 15 -237 25
rect -329 14 -237 15
rect -329 -2 -262 14
rect -329 -52 -312 -2
rect -268 -3 -262 -2
rect -245 -3 -237 14
rect -268 -11 -237 -3
rect -181 19 -163 53
rect -122 19 -105 53
rect -181 2 -105 19
rect -181 -52 -163 2
rect -122 -52 -105 2
rect -87 16 -57 24
rect -87 -1 -81 16
rect -64 -1 -57 16
rect -87 -9 -57 -1
rect -35 -52 -18 53
rect -741 -60 -707 -52
rect -741 -77 -733 -60
rect -716 -77 -707 -60
rect -741 -82 -707 -77
rect -673 -57 -640 -52
rect -673 -74 -666 -57
rect -649 -74 -640 -57
rect -673 -82 -640 -74
rect -568 -57 -535 -52
rect -568 -74 -560 -57
rect -543 -74 -535 -57
rect -568 -82 -535 -74
rect -497 -58 -464 -52
rect -497 -75 -489 -58
rect -472 -75 -464 -58
rect -497 -82 -464 -75
rect -403 -60 -369 -52
rect -403 -77 -395 -60
rect -378 -77 -369 -60
rect -403 -82 -369 -77
rect -335 -57 -302 -52
rect -335 -74 -328 -57
rect -311 -74 -302 -57
rect -335 -82 -302 -74
rect -256 -59 -223 -52
rect -256 -76 -248 -59
rect -231 -76 -223 -59
rect -256 -82 -223 -76
rect -189 -60 -155 -52
rect -189 -77 -180 -60
rect -163 -77 -155 -60
rect -189 -82 -155 -77
rect -122 -58 -89 -52
rect -122 -75 -114 -58
rect -97 -75 -89 -58
rect -122 -82 -89 -75
rect -51 -58 -18 -52
rect -51 -75 -43 -58
rect -26 -75 -18 -58
rect -51 -82 -18 -75
rect 20 91 51 99
rect 20 61 27 91
rect 45 61 51 91
rect 20 53 51 61
rect 93 91 124 99
rect 93 61 100 91
rect 118 61 124 91
rect 93 53 124 61
rect 160 91 194 99
rect 160 61 168 91
rect 186 61 194 91
rect 160 53 194 61
rect 230 91 264 99
rect 230 61 238 91
rect 256 61 264 91
rect 230 53 264 61
rect 299 91 333 99
rect 299 61 308 91
rect 326 61 333 91
rect 299 53 333 61
rect 369 91 403 99
rect 369 61 378 91
rect 396 61 403 91
rect 369 53 403 61
rect 439 91 470 99
rect 439 61 445 91
rect 463 61 470 91
rect 439 53 470 61
rect 512 91 543 99
rect 512 61 518 91
rect 536 61 543 91
rect 512 53 543 61
rect 20 -52 37 53
rect 57 23 87 31
rect 57 6 63 23
rect 80 6 87 23
rect 57 -2 87 6
rect 107 16 124 53
rect 146 16 181 22
rect 107 -1 155 16
rect 172 -1 181 16
rect 107 -52 124 -1
rect 146 -9 181 -1
rect 236 16 253 53
rect 285 16 320 23
rect 236 -1 294 16
rect 311 -1 320 16
rect 236 -52 253 -1
rect 285 -8 320 -1
rect 375 17 392 53
rect 439 17 456 53
rect 375 0 456 17
rect 375 -52 392 0
rect 439 -52 456 0
rect 477 -10 507 -2
rect 477 -27 483 -10
rect 500 -27 507 -10
rect 477 -35 507 -27
rect 526 -52 543 53
rect 20 -57 52 -52
rect 20 -74 27 -57
rect 44 -74 52 -57
rect 20 -82 52 -74
rect 92 -59 124 -52
rect 92 -76 100 -59
rect 117 -76 124 -59
rect 92 -82 124 -76
rect 162 -60 196 -52
rect 162 -77 170 -60
rect 187 -77 196 -60
rect 162 -82 196 -77
rect 230 -57 263 -52
rect 230 -74 237 -57
rect 254 -74 263 -57
rect 230 -82 263 -74
rect 301 -60 335 -52
rect 301 -77 309 -60
rect 326 -77 335 -60
rect 301 -82 335 -77
rect 369 -57 402 -52
rect 369 -74 376 -57
rect 393 -74 402 -57
rect 369 -82 402 -74
rect 439 -57 471 -52
rect 439 -74 446 -57
rect 463 -74 471 -57
rect 439 -82 471 -74
rect 511 -58 543 -52
rect 511 -75 519 -58
rect 536 -75 543 -58
rect 511 -82 543 -75
rect -735 -150 -718 -82
rect -481 -96 -464 -82
rect -397 -150 -380 -82
rect -249 -150 -232 -82
rect -35 -93 -18 -82
rect -35 -112 -18 -110
rect 107 -92 124 -82
rect 107 -111 124 -109
rect 168 -150 185 -82
rect 307 -150 324 -82
rect 526 -93 543 -82
rect 526 -114 543 -111
rect -744 -167 -735 -150
rect -718 -167 -710 -150
rect -693 -167 -397 -150
rect -380 -167 -374 -150
rect -357 -167 -278 -150
rect -261 -167 -249 -150
rect -232 -167 168 -150
rect 185 -167 196 -150
rect 213 -167 273 -150
rect 290 -167 307 -150
rect 324 -167 341 -150
<< viali >>
rect -735 191 -718 208
rect -397 191 -380 208
rect -252 191 -235 208
rect 168 191 185 208
rect 307 191 324 208
rect -209 138 -192 155
rect 20 135 37 152
rect -787 26 -770 43
rect -606 24 -589 41
rect -644 -28 -627 -11
rect -525 -28 -508 -11
rect -81 -1 -64 16
rect 63 6 80 23
rect 483 -27 500 -10
rect -481 -113 -464 -96
rect -35 -110 -18 -93
rect 107 -109 124 -92
rect 526 -111 543 -93
rect -735 -167 -718 -150
rect -397 -167 -380 -150
rect -249 -167 -232 -150
rect 168 -167 185 -150
rect 307 -167 324 -150
<< metal1 >>
rect -755 208 364 217
rect -755 191 -735 208
rect -718 191 -397 208
rect -380 191 -252 208
rect -235 191 168 208
rect 185 191 307 208
rect 324 191 364 208
rect -755 180 364 191
rect -755 179 -632 180
rect -221 155 43 163
rect -221 138 -209 155
rect -192 152 43 155
rect -192 138 20 152
rect -221 135 20 138
rect 37 135 43 152
rect -221 129 43 135
rect -793 43 -583 48
rect -793 26 -787 43
rect -770 41 -583 43
rect -770 26 -606 41
rect -793 24 -606 26
rect -589 24 -583 41
rect -793 17 -583 24
rect -90 16 -53 24
rect -90 -1 -81 16
rect -64 -1 -53 16
rect 54 23 91 26
rect 54 6 63 23
rect 80 6 91 23
rect 54 -1 91 6
rect -650 -10 508 -1
rect -650 -11 483 -10
rect -650 -28 -644 -11
rect -627 -28 -525 -11
rect -508 -27 483 -11
rect 500 -27 508 -10
rect -508 -28 508 -27
rect -650 -35 508 -28
rect -489 -93 -9 -88
rect -489 -96 -35 -93
rect -489 -113 -481 -96
rect -464 -110 -35 -96
rect -18 -110 -9 -93
rect -464 -113 -9 -110
rect -489 -116 -9 -113
rect 101 -92 549 -86
rect 101 -109 107 -92
rect 124 -93 549 -92
rect 124 -109 526 -93
rect 101 -111 526 -109
rect 543 -111 549 -93
rect 101 -114 549 -111
rect -749 -150 341 -144
rect -749 -167 -735 -150
rect -718 -167 -397 -150
rect -380 -167 -249 -150
rect -232 -167 168 -150
rect 185 -167 307 -150
rect 324 -167 341 -150
rect -749 -175 341 -167
<< labels >>
flabel locali -667 -28 -649 -11 0 FreeSans 72 0 0 0 clkbar
flabel locali -304 -2 -286 15 0 FreeSans 80 0 0 0 2
flabel locali -155 2 -138 19 0 FreeSans 80 0 0 0 3
flabel locali 107 -1 124 16 0 FreeSans 80 0 0 0 4
flabel locali 401 0 420 17 0 FreeSans 80 0 0 0 5
flabel metal1 -611 192 -554 207 0 FreeSans 152 0 0 0 vdd
flabel metal1 -661 -166 -589 -150 0 FreeSans 152 0 0 0 gnd
flabel locali -808 27 -794 42 0 FreeSans 120 0 0 0 din
flabel locali 236 -1 266 16 0 FreeSans 120 0 0 0 Q
flabel locali -777 -24 -755 -9 0 FreeSans 120 0 0 0 clk
flabel locali -464 -1 -434 16 0 FreeSans 120 0 0 0 1
<< end >>
