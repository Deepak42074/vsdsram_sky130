*Description of Tristate Buffer
.param temp=27
.param supl = 1.8V

*Including sky130 devoce models
.lib "sky130_fd_pr/models/sky130.lib.spice" tt

Vdd vdd 0 {supl}

* transistors
*inverter

XM1 inb in vdd vdd sky130_fd_pr__pfet_01v8 w=.42 l=.15 m=1
XM2 inb in 0 0 sky130_fd_pr__nfet_01v8 w=.42 l=.15 m=1

XM3 out1 inb vdd vdd sky130_fd_pr__pfet_01v8 w=.42 l=.15 m=1
XM4 out1 inb 0 0 sky130_fd_pr__nfet_01v8 w=.42 l=.15 m=1

XM5 out enb out1 vdd sky130_fd_pr__pfet_01v8 w=.55 l=.15 m=1
XM6 out en out1 0  sky130_fd_pr__nfet_01v8 w=.55 l=.15 m=1

*Pull down ckt for Transmission gate is disabled case
XM7 out enb 0 0  sky130_fd_pr__nfet_01v8 w=.55 l=.15 m=1

* Sources
Vin in 0 pulse(0 1.8 0 60ps 60ps 0.5ns 1ns)
Ven en 0 pulse(0 1.8 0 60ps 60ps 2ns 4ns)
Venb enb 0 pulse(1.8 0 0 60ps 60ps 2ns 4ns)

.tran 0.01p 10ns

.control
run

plot en+6 enb+4 in+2 out
.endc
.end




 


